module COUNT24 (RESET, CLK, LED7seg, SEL_DOWN, SA, BTN1, BTN2, BTN3, CS_COLOR1, CS_COLOR2, CS_COLOR3);
input RESET, CLK, SEL_DOWN, BTN1, BTN2, BTN3;
output [7:0] LED7seg;
output [3:0] SA;
output [3:0] CS_COLOR1;
output [2:0] CS_COLOR2, CS_COLOR3;


parameter SETTIME1_MAX = 125000000; // 125MHz


wire ENABLE, ENABLE_kHz, EN05, BAP_BTN1, BAP_BTN2, BAP_BTN3, ALARM_ON, ALARM_STATE;
wire [6:0] SETUP_TIME, SETUP_ALARM;
wire [4:0] SEL_MODE;
wire [3:0] COUNT_10, COUNT_10m, COUNT_10h, ACOUNT_10m, ACOUNT_10h;
wire [2:0] COUNT_6, COUNT_6m, ACOUNT_6m;
wire [1:0] COUNT_2h, ACOUNT_2h, CURRENT_STATE_TIME;

wire [3:0] LED_COUNT;
wire [3:0] L1, L2, L3, L4;
wire CARRY59;
wire CARRY5959;

secCOUNT i0(.RESET(RESET), .CLK(CLK), .ENABLE(ENABLE), .ENABLE_kHz(ENABLE_kHz), .EN05(EN05));
SETUP_SW i1(.CLK(CLK), .ENABLE_kHz(ENABLE_kHz), .BTN(BTN1), .BAP_BTN(BAP_BTN1));
SETUP_SW i2(.CLK(CLK), .ENABLE_kHz(ENABLE_kHz), .BTN(BTN2), .BAP_BTN(BAP_BTN2));
SETUP_SW i3(.CLK(CLK), .ENABLE_kHz(ENABLE_kHz), .BTN(BTN3), .BAP_BTN(BAP_BTN3));
SEQ_SELMODE i10(.RESET(RESET), .CLK(CLK), .BAP_BTN1(BAP_BTN1), .CURRENT_STATE_TIME(SEL_MODE));
SEQ_SET_TIME i11(.RESET(RESET), .CLK(CLK), .BAP_BTN2(BAP_BTN2), .CURRENT_STATE_TIME(SETUP_TIME), .SEL_MODE0(SEL_MODE[0]));
SEQUENCER i12(.RESET(RESET), .CLK(CLK), .BAP_BTN3(BAP_BTN3), .CURRENT_STATE_TIME(CURRENT_STATE_TIME), .SEL_MODE1(SEL_MODE[1]));
//new
SEQ_SET_ALARM i13(.RESET(RESET), .CLK(CLK), .BAP_BTN2(BAP_BTN2), .CURRENT_STATE_TIME(SETUP_ALARM), .SEL_MODE2(SEL_MODE[2]));
SEQ_ALARM_USE i14(.RESET(RESET), .CLK(CLK), .BAP_BTN3(BAP_BTN3), .ALARM_ON(ALARM_ON), .SEL_MODE2(SEL_MODE[2]), .SETUP_ALARM0(SETUP_ALARM[0]));
//

CNT60 i20(.RESET(RESET), .CLK(CLK), .SEL_DOWN(SEL_DOWN), .COUNT_10(COUNT_10), .COUNT_6(COUNT_6), 
         .ENABLE(ENABLE), .CIN({1'b1}), .COUT(CARRY59), .BASE(SETUP_TIME[0]), 
         .SETTIME1(SETUP_TIME[6]), .SETTIME10(SETUP_TIME[5]), .BAP_BTN3(BAP_BTN3));
CNT60 i21(.RESET(RESET), .CLK(CLK), .SEL_DOWN(SEL_DOWN), .COUNT_10(COUNT_10m), .COUNT_6(COUNT_6m), 
         .ENABLE(ENABLE), .CIN(CARRY59), .COUT(CARRY5959), .BASE(SETUP_TIME[0]),
         .SETTIME1(SETUP_TIME[4]), .SETTIME10(SETUP_TIME[3]), .BAP_BTN3(BAP_BTN3));
CNT24 i22(.RESET(RESET), .CLK(CLK), .SEL_DOWN(SEL_DOWN), .COUNT_10(COUNT_10h), .COUNT_2(COUNT_2h), 
         .ENABLE(ENABLE), .CIN(CARRY5959), .COUT(), .BASE(SETUP_TIME[0]),
         .SETTIME1(SETUP_TIME[2]), .SETTIME10(SETUP_TIME[1]), .BAP_BTN3(BAP_BTN3));
//new
CNT60_ALARM i23(.RESET(RESET), .CLK(CLK), .SEL_DOWN(SEL_DOWN), .COUNT_10(ACOUNT_10m), .COUNT_6(ACOUNT_6m), 
                .SETTIME1(SETUP_ALARM[4]), .SETTIME10(SETUP_ALARM[3]), .BAP_BTN3(BAP_BTN3));
CNT24_ALARM i24(.RESET(RESET), .CLK(CLK), .SEL_DOWN(SEL_DOWN), .COUNT_10(ACOUNT_10h), .COUNT_2(ACOUNT_2h), 
                .SETTIME1(SETUP_ALARM[2]), .SETTIME10(SETUP_ALARM[1]), .BAP_BTN3(BAP_BTN3));
//

DE_SELECTER i30(.RESET(RESET), .CLK(CLK),
                .SEL(CURRENT_STATE_TIME), .L1(L1), .L2(L2), .L3(L3), .L4(L4),
                .COUNT_10(COUNT_10), .COUNT_10m(COUNT_10m), .COUNT_10h(COUNT_10h), .COUNT_6(COUNT_6), .COUNT_6m(COUNT_6m), .COUNT_2h(COUNT_2h),
                .EN05(EN05), .SEL_MODE(SEL_MODE), .SETUP_TIME(SETUP_TIME),
                .ACOUNT_10m(ACOUNT_10m), .ACOUNT_10h(ACOUNT_10h), .ACOUNT_6m(ACOUNT_6m), .ACOUNT_2h(ACOUNT_2h),
                .BAP_BTN1(BAP_BTN1), .SETUP_ALARM(SETUP_ALARM[4:0]), .ALARM_STATE(ALARM_STATE), .ALARM_ON(ALARM_ON)); 

DCOUNT  i31(.RESET(RESET), .CLK(CLK), .ENABLE_kHz(ENABLE_kHz), .L1(L1), .L2(L2),
            .L3(L3), .L4(L4), .SA(SA), .L(LED_COUNT));
DECODER i32(.LED_COUNT(LED_COUNT), .LED7seg(LED7seg));

LED_COLOR1 i40(.SETUP_TIME(SETUP_TIME), .CURRENT_STATE_LED(CS_COLOR1));
LED_COLOR2 i41(.SEL_MODE(SEL_MODE), .CURRENT_STATE_COLOR(CS_COLOR2));
LED_COLOR3 i42(.ALARM_STATE(ALARM_STATE), .CURRENT_STATE_COLOR(CS_COLOR3));

endmodule